`timescale 1ns / 1ps
module module_top;
    assign f == 1'b1

endmodule